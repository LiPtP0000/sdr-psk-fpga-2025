// Module: PSK_Signal_Extend
// =========================
// This module extends the PSK signal to a wider width. (Actually not used now, when I_WIDTH == Q_WIDTH).
// It also allows the selection of I or Q stream for later processing.
//
// Author: LiPtP
// Date: 2025/12/18

`timescale 1ns / 1ps

module PSK_Signal_Extend #(
    parameter I_WIDTH    = 12,
    parameter O_WIDTH    = 16,
    parameter USE_I_STRM = 1 // 1 for I stream, 0 for Q stream
) (
    input                           clk,
    input  signed     [I_WIDTH-1:0] DAC_I,
    input  signed     [I_WIDTH-1:0] DAC_Q,
    input                           is_bpsk,
    output reg signed [O_WIDTH-1:0] PSK_signal,
    output reg                      is_bpsk_out
);
    reg signed [O_WIDTH-1:0] PSK_signal_d;
    reg                      is_bpsk_out_d;

    // assign LSB to zeros
    generate
        if (USE_I_STRM) begin
            always @(posedge clk) begin
                PSK_signal_d <= {DAC_I, {O_WIDTH - I_WIDTH{1'b0}}};
            end
        end else begin
            always @(posedge clk) begin
                PSK_signal_d <= {DAC_Q, {O_WIDTH - I_WIDTH{1'b0}}};
            end
        end
    endgenerate

    always @(posedge clk) begin
        is_bpsk_out_d <= is_bpsk;

        PSK_signal    <= PSK_signal_d;
        is_bpsk_out   <= is_bpsk_out_d;
    end
endmodule
