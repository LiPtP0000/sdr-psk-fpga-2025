module Rx_wrapper (
    input         clk_1M024,
    input         clk_2M048,
    input         clk_16M384,
    input         clk_32M768,
    input  [11:0] ADC_I,
    input  [11:0] ADC_Q,
    input         rst_16M384,
    input         rst_32M768,
    input  [ 3:0] MODE_CTRL,
    input  [ 3:0] FEEDBACK_SHIFT,
    input  [ 3:0] GARDNER_SHIFT,
    input  [15:0] RX_SD_THRESHOLD,
    input  [ 7:0] RX_SD_WINDOW,
    input  [ 7:0] RX_PD_WINDOW,
    input  [ 7:0] RX_BD_WINDOW,
    output        BPSK_raw,
    output [ 1:0] QPSK_raw,
    output [15:0] I_16M,
    output [15:0] Q_16M,
    output [11:0] NCO_cos,
    output [15:0] I_1M,
    output [15:0] Q_1M,
    output        clk_1M_out,
    output [ 1:0] QPSK,
    output        BPSK,
    output        Rx_1bit,
    output [ 7:0] data_tdata,
    output        data_tvalid,
    output        data_tlast,
    output        data_tuser,
    output [15:0] error_tdata,
    output [15:0] feedback_tdata,
    output        Rx_valid,
    output [15:0] gardner_error,
    output [15:0] gardner_increment
);

// 
endmodule
